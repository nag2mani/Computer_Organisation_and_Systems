//This is for XOR logic.
module xor_logic(a, b, c);
input a,b;
output c;
assign c = a ^ b;
endmodule
