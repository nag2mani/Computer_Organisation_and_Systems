//This is for and logic.

module and_logic(a, b, c);
input a, b;
output c;
assign c = a & b;
endmodule
