//This is for or logic.
module or_logic(a, b, c);
input a, b;
output c;
assign c = a | b;
endmodule
