//This is for not logic.
module not_logic(a, b); //Here a is input and b is output.
input a;
output b;
assign b = ~a;
endmodule
